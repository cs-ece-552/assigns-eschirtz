/*
    CS/ECE 552 Spring '19
    Homework #3, Problem 2

    1 input NOT
*/
module not1 (in1,out);
    input in1;
    output out;
    assign out = ~in1;
endmodule