s/*
   CS/ECE 552, Spring '19
   Homework #6, Problem #1
  
   This module determines all of the control logic for the processor.
*/
module control (/*AUTOARG*/
                // Outputs
                err, 
                RegDst,
                SESel,
                RegWrite,
                DMemWrite,
                DMemEn,
                ALUSrc2,
                PCSrc,
                MemToReg,
                DMemDump,
                Jump,
                // Inputs
                OpCode,
                Funct
                );

   // inputs
   input [4:0]  OpCode;
   input [1:0]  Funct;
   
   // outputs
   output       err;
   output       RegDst, RegWrite, DMemWrite, DMemEn, ALUSrc2, PCSrc, 
                MemToReg, DMemDump, Jump;
   output [1:0] RegDst;
   output [2:0] SESel;

   /* YOUR CODE HERE */
   
endmodule
